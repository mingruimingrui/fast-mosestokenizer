#single upper case letter are usually initials
A
B
C
D
E
F
G
H
I
J
K
L
M
N
O
P
Q
R
S
T
U
V
W
X
Y
Z
Å
Ä
Ö
#misc abbreviations
#If all words in text are in small case, then tex, mao, tom, maj, may be confused with names, and iaf, etc with named entities.
AB
VG
dvs
d.v.s
d. v. s
etc
from
fr.o.m
fr. o. m
iaf
i.a.f
i. a. f
jfr
kl
kr
mao
m.a.o
m. a. o
mfl
m.fl
m. fl
mm
m.m
m. m.
osv
o.s.v
o. s. v
pga
p.g.a
p. g. a
tex
t.ex
t. ex
#tom. is risky, as tom is a word, and can be at end of sentence. One recent text has 9 tom., and 52 tom not at end of sentence.
tom
t.o.m
t. o. m
vs
adv
jur
kand
mag
fil
lic
prop
d
f
s
mha
m.h.a
m. h. a
vol
#months
jan
feb
mar
apr
#maj is a full word
jun
jul
aug
sep
okt
nov
dec
